module delay_clap(
  input clk_1,
  input rst_n,
  input signal_1,
  input clk_2,
  output signal_2
);
